module top_module ( input a,b, output out);
  assign = !(a^b);
endmodule
